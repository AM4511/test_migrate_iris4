/****************************************************************************
 * core_pkg.sv
 ****************************************************************************/

/**
 * Package: core_pkg
 *
 * TODO: Add package documentation
 */
package core_pkg;
	// this is a forward type definition (For the `include section below)
	typedef class Cstatus;

	`include "Cstatus.svh"

endpackage