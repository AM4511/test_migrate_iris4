/****************************************************************************
 * registerfile_pkg.sv
 ****************************************************************************/

/**
 * Package: registerfile_pkg
 * 
 * TODO: Add package documentation
 */
package registerfile_pkg;
	
	typedef class Cnode;
//	typedef class Cregisterfile;
//	typedef class Csection;
//	typedef class Cexternal;
//	typedef class Cregister;
//	typedef class Cfield;


	`include "Cnode.svh"
//	`include "Cregisterfile.svh"
//	`include "Csection.svh"
//	`include "Cexternal.svh"
//	`include "Cregister.svh"
//	`include "Cfield.svh"

endpackage


