/****************************************************************************
 * fdkide_pkg.sv
 ****************************************************************************/

/**
 * Package: fdkide_pkg
 * 
 * TODO: Add package documentation
 */
package athena_pkg;

	typedef class Cathena;
	
	`include "Cathena.svh"

	
endpackage


