/****************************************************************************
 * dmawr2tlp_pkg.sv
 ****************************************************************************/

/**
 * Package: dmawr2tlp_pkg
 *
 * TODO: Add package documentation
 */

package dmawr2tlp_pkg;
	import core_pkg::*;
	import driver_pkg::*;

	typedef class Cscoreboard_dmawr2tlp;
	
	`include "Cscoreboard_dmawr2tlp.svh"

endpackage : dmawr2tlp_pkg








