/****************************************************************************
 * test_pkg.sv
 ****************************************************************************/

/**
 * Package: tests_pkg
 *
 * TODO: Add package documentation
 */
package tests_pkg;
    
  `include "test0001.svh"
  `include "test0002.svh"
  `include "test0003.svh"
  `include "test0004.svh"
  `include "test0005.svh"
  `include "test0006.svh"
  `include "test0007.svh"
  `include "test0008.svh"
  `include "test0009.svh"
  `include "test0010.svh"
  `include "test0020.svh"
  `include "test0021.svh"
  `include "test0022.svh"
  `include "test0023.svh"  
  `include "test0024.svh"   
  `include "test0025.svh"   
  
  typedef class Test0001;
  typedef class Test0002;  
  typedef class Test0003;    
  typedef class Test0004;   
  typedef class Test0005; 
  typedef class Test0006;   
  typedef class Test0007;
  typedef class Test0008;
  typedef class Test0009;
  typedef class Test0010;
  typedef class Test0020;
  typedef class Test0021;
  typedef class Test0022;    
  typedef class Test0023;     
  typedef class Test0024; 
  typedef class Test0025;     

endpackage
