/****************************************************************************
 * xgs_pkg.sv
 ****************************************************************************/

/**
 * Package: xgs_pkg
 * 
 * TODO: Add package documentation
 */
package xgs_pkg;
	typedef class Cxgs_sensor;
	typedef class Cxgs12M;

	`include "Cxgs_sensor.svh"
    `include "Cxgs12M.svh"
endpackage


