/****************************************************************************
 * image_pkg.sv
 ****************************************************************************/

/**
 * Package: image_pkg
 *
 * TODO: Add package documentation
 */

package image_pkg;

	typedef class Cimage;
	
	`include "Cimage.svh"
endpackage








