hispi_phy_altera_inst : hispi_phy_altera PORT MAP (
		pll_areset	 => pll_areset_sig,
		rx_in	 => rx_in_sig,
		rx_inclock	 => rx_inclock_sig,
		rx_locked	 => rx_locked_sig,
		rx_out	 => rx_out_sig,
		rx_outclock	 => rx_outclock_sig
	);
