/****************************************************************************
 * Csensor.svh
 ****************************************************************************/

/**
 * Class: Csensor
 * 
 * TODO: Add class documentation
 */
class Csensor;

	function new();

	endfunction


endclass


