/****************************************************************************
 * fpga_cfg_pkg.sv
 ****************************************************************************/

/**
 * Package: fpga_cfg_pkg
 *
 * TODO: Add package documentation
 */
package fpga_cfg_pkg;
    
parameter COLOR = 0;
    
endpackage
