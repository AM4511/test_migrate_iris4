/****************************************************************************
 * driver_pkg.sv
 ****************************************************************************/

/**
 * Package: driver_pkg
 *
 * TODO: Add package documentation
 */
package driver_pkg;

	`include "Cdriver_axil.svh"

	typedef class Cdriver_axil;



endpackage


