/****************************************************************************
 * img_testpack.sv
 ****************************************************************************/

/**
 * Package: tests_pkg
 *
 * TODO: Add package documentation
 */
package tests_pkg;
	typedef class Ctest0000;

//	typedef class Ctest0001;
//	typedef class Ctest0002;
//	typedef class Ctest0003;
//	typedef class Ctest0004;
//	typedef class Ctest0005;
//	typedef class Ctest0006;
//	typedef class Ctest0010;
//	typedef class Ctest0011;
	typedef class Ctest0100;
	typedef class Ctest0101;
	typedef class Ctest0110;
	typedef class Ctest0200;
	typedef class Ctest0300;
	typedef class Ctest0400;
	typedef class Ctest0500;
	typedef class CtestManager;

//	`include "Ctest0001.svh"
//	`include "Ctest0002.svh"
//	`include "Ctest0003.svh"
//	`include "Ctest0004.svh"
//	`include "Ctest0005.svh"
//	`include "Ctest0006.svh"
//	`include "Ctest0010.svh"
//	`include "Ctest0011.svh"
	`include "registerfile/Ctest0000.svh"
	`include "timers/Ctest0400.svh"
	`include "io/Ctest0500.svh"
	`include "Ctest0100.svh"
	`include "Ctest0101.svh"
	`include "Ctest0110.svh"
	`include "Ctest0200.svh"
	`include "Ctest0300.svh"
	`include "CtestManager.svh"

endpackage


