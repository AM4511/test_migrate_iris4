library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


package hispi_pack is
  -- constant HISPI_PIXEL_SIZE    : integer := 20;
  -- constant MAX_PIXELS_PER_LINE : integer := 1280;
  -- constant MAX_LINES_PER_FRAME : integer := 960;



end package hispi_pack;

package body hispi_pack is



end package body hispi_pack;
