/****************************************************************************
 * Csection.svh
 ****************************************************************************/

/**
 * Class: Csection
 * 
 * TODO: Add class documentation
 */
class Csection extends Cnode;
	
	function new(Cnode parent = null, longint offset=0);
		super.new(parent, offset);
	endfunction


endclass


