/****************************************************************************
 * xgs_athena_pkg.sv
 ****************************************************************************/

/**
 * Package: xgs_athena_pkg
 *
 * TODO: Add package documentation
 */

package xgs_athena_pkg;
	import core_pkg::*;
	import driver_pkg::*;
	
	typedef class CImage;
	`include "Cimage.sv"
	
	typedef class Cscoreboard;
	`include "Cscoreboard.svh"


	
endpackage : xgs_athena_pkg








